`timescale 1ns / 1ps
//////////////////////////////////////////////////////////////////////////////////
// Company: 
// Engineer: 
// 
// Create Date:    16:28:16 08/27/2017 
// Design Name: 
// Module Name:    reduction_table_q60bit 
// Project Name: 
// Target Devices: 
// Tool versions: 
// Description: 
//
// Dependencies: 
//
// Revision: 
// Revision 0.01 - File Created
// Additional Comments: 
//
//////////////////////////////////////////////////////////////////////////////////
module reduction_table_q1068564481(i, table_out);
input [5:0] i;
output [29:0] table_out;
assign table_out = 
   (i==6'd0) ? 30'd0 :
   (i==6'd1) ? 30'd5177343 :
   (i==6'd2) ? 30'd10354686 :
   (i==6'd3) ? 30'd15532029 :
   (i==6'd4) ? 30'd20709372 :
   (i==6'd5) ? 30'd25886715 :
   (i==6'd6) ? 30'd31064058 :
   (i==6'd7) ? 30'd36241401 :
   (i==6'd8) ? 30'd41418744 :
   (i==6'd9) ? 30'd46596087 :
   (i==6'd10) ? 30'd51773430 :
   (i==6'd11) ? 30'd56950773 :
   (i==6'd12) ? 30'd62128116 :
   (i==6'd13) ? 30'd67305459 :
   (i==6'd14) ? 30'd72482802 :
   (i==6'd15) ? 30'd77660145 :
   (i==6'd16) ? 30'd82837488 :
   (i==6'd17) ? 30'd88014831 :
   (i==6'd18) ? 30'd93192174 :
   (i==6'd19) ? 30'd98369517 :
   (i==6'd20) ? 30'd103546860 :
   (i==6'd21) ? 30'd108724203 :
   (i==6'd22) ? 30'd113901546 :
   (i==6'd23) ? 30'd119078889 :
   (i==6'd24) ? 30'd124256232 :
   (i==6'd25) ? 30'd129433575 :
   (i==6'd26) ? 30'd134610918 :
   (i==6'd27) ? 30'd139788261 :
   (i==6'd28) ? 30'd144965604 :
   (i==6'd29) ? 30'd150142947 :
   (i==6'd30) ? 30'd155320290 :
   (i==6'd31) ? 30'd160497633 :
   (i==6'd32) ? 30'd165674976 :
   (i==6'd33) ? 30'd170852319 :
   (i==6'd34) ? 30'd176029662 :
   (i==6'd35) ? 30'd181207005 :
   (i==6'd36) ? 30'd186384348 :
   (i==6'd37) ? 30'd191561691 :
   (i==6'd38) ? 30'd196739034 :
   (i==6'd39) ? 30'd201916377 :
   (i==6'd40) ? 30'd207093720 :
   (i==6'd41) ? 30'd212271063 :
   (i==6'd42) ? 30'd217448406 :
   (i==6'd43) ? 30'd222625749 :
   (i==6'd44) ? 30'd227803092 :
   (i==6'd45) ? 30'd232980435 :
   (i==6'd46) ? 30'd238157778 :
   (i==6'd47) ? 30'd243335121 :
   (i==6'd48) ? 30'd248512464 :
   (i==6'd49) ? 30'd253689807 :
   (i==6'd50) ? 30'd258867150 :
   (i==6'd51) ? 30'd264044493 :
   (i==6'd52) ? 30'd269221836 :
   (i==6'd53) ? 30'd274399179 :
   (i==6'd54) ? 30'd279576522 :
   (i==6'd55) ? 30'd284753865 :
   (i==6'd56) ? 30'd289931208 :
   (i==6'd57) ? 30'd295108551 :
   (i==6'd58) ? 30'd300285894 :
   (i==6'd59) ? 30'd305463237 :
   (i==6'd60) ? 30'd310640580 :
   (i==6'd61) ? 30'd315817923 :
   (i==6'd62) ? 30'd320995266 :
   30'd326172609;

endmodule


module reduction_table_q1069219841(i, table_out);
input [5:0] i;
output [29:0] table_out;
assign table_out = 
   (i==6'd0) ? 30'd0 :
   (i==6'd1) ? 30'd4521983 :
   (i==6'd2) ? 30'd9043966 :
   (i==6'd3) ? 30'd13565949 :
   (i==6'd4) ? 30'd18087932 :
   (i==6'd5) ? 30'd22609915 :
   (i==6'd6) ? 30'd27131898 :
   (i==6'd7) ? 30'd31653881 :
   (i==6'd8) ? 30'd36175864 :
   (i==6'd9) ? 30'd40697847 :
   (i==6'd10) ? 30'd45219830 :
   (i==6'd11) ? 30'd49741813 :
   (i==6'd12) ? 30'd54263796 :
   (i==6'd13) ? 30'd58785779 :
   (i==6'd14) ? 30'd63307762 :
   (i==6'd15) ? 30'd67829745 :
   (i==6'd16) ? 30'd72351728 :
   (i==6'd17) ? 30'd76873711 :
   (i==6'd18) ? 30'd81395694 :
   (i==6'd19) ? 30'd85917677 :
   (i==6'd20) ? 30'd90439660 :
   (i==6'd21) ? 30'd94961643 :
   (i==6'd22) ? 30'd99483626 :
   (i==6'd23) ? 30'd104005609 :
   (i==6'd24) ? 30'd108527592 :
   (i==6'd25) ? 30'd113049575 :
   (i==6'd26) ? 30'd117571558 :
   (i==6'd27) ? 30'd122093541 :
   (i==6'd28) ? 30'd126615524 :
   (i==6'd29) ? 30'd131137507 :
   (i==6'd30) ? 30'd135659490 :
   (i==6'd31) ? 30'd140181473 :
   (i==6'd32) ? 30'd144703456 :
   (i==6'd33) ? 30'd149225439 :
   (i==6'd34) ? 30'd153747422 :
   (i==6'd35) ? 30'd158269405 :
   (i==6'd36) ? 30'd162791388 :
   (i==6'd37) ? 30'd167313371 :
   (i==6'd38) ? 30'd171835354 :
   (i==6'd39) ? 30'd176357337 :
   (i==6'd40) ? 30'd180879320 :
   (i==6'd41) ? 30'd185401303 :
   (i==6'd42) ? 30'd189923286 :
   (i==6'd43) ? 30'd194445269 :
   (i==6'd44) ? 30'd198967252 :
   (i==6'd45) ? 30'd203489235 :
   (i==6'd46) ? 30'd208011218 :
   (i==6'd47) ? 30'd212533201 :
   (i==6'd48) ? 30'd217055184 :
   (i==6'd49) ? 30'd221577167 :
   (i==6'd50) ? 30'd226099150 :
   (i==6'd51) ? 30'd230621133 :
   (i==6'd52) ? 30'd235143116 :
   (i==6'd53) ? 30'd239665099 :
   (i==6'd54) ? 30'd244187082 :
   (i==6'd55) ? 30'd248709065 :
   (i==6'd56) ? 30'd253231048 :
   (i==6'd57) ? 30'd257753031 :
   (i==6'd58) ? 30'd262275014 :
   (i==6'd59) ? 30'd266796997 :
   (i==6'd60) ? 30'd271318980 :
   (i==6'd61) ? 30'd275840963 :
   (i==6'd62) ? 30'd280362946 :
   30'd284884929;

endmodule


module reduction_table_q1070727169(i, table_out);
input [5:0] i;
output [29:0] table_out;
assign table_out = 
   (i==6'd0) ? 30'd0 :
   (i==6'd1) ? 30'd3014655 :
   (i==6'd2) ? 30'd6029310 :
   (i==6'd3) ? 30'd9043965 :
   (i==6'd4) ? 30'd12058620 :
   (i==6'd5) ? 30'd15073275 :
   (i==6'd6) ? 30'd18087930 :
   (i==6'd7) ? 30'd21102585 :
   (i==6'd8) ? 30'd24117240 :
   (i==6'd9) ? 30'd27131895 :
   (i==6'd10) ? 30'd30146550 :
   (i==6'd11) ? 30'd33161205 :
   (i==6'd12) ? 30'd36175860 :
   (i==6'd13) ? 30'd39190515 :
   (i==6'd14) ? 30'd42205170 :
   (i==6'd15) ? 30'd45219825 :
   (i==6'd16) ? 30'd48234480 :
   (i==6'd17) ? 30'd51249135 :
   (i==6'd18) ? 30'd54263790 :
   (i==6'd19) ? 30'd57278445 :
   (i==6'd20) ? 30'd60293100 :
   (i==6'd21) ? 30'd63307755 :
   (i==6'd22) ? 30'd66322410 :
   (i==6'd23) ? 30'd69337065 :
   (i==6'd24) ? 30'd72351720 :
   (i==6'd25) ? 30'd75366375 :
   (i==6'd26) ? 30'd78381030 :
   (i==6'd27) ? 30'd81395685 :
   (i==6'd28) ? 30'd84410340 :
   (i==6'd29) ? 30'd87424995 :
   (i==6'd30) ? 30'd90439650 :
   (i==6'd31) ? 30'd93454305 :
   (i==6'd32) ? 30'd96468960 :
   (i==6'd33) ? 30'd99483615 :
   (i==6'd34) ? 30'd102498270 :
   (i==6'd35) ? 30'd105512925 :
   (i==6'd36) ? 30'd108527580 :
   (i==6'd37) ? 30'd111542235 :
   (i==6'd38) ? 30'd114556890 :
   (i==6'd39) ? 30'd117571545 :
   (i==6'd40) ? 30'd120586200 :
   (i==6'd41) ? 30'd123600855 :
   (i==6'd42) ? 30'd126615510 :
   (i==6'd43) ? 30'd129630165 :
   (i==6'd44) ? 30'd132644820 :
   (i==6'd45) ? 30'd135659475 :
   (i==6'd46) ? 30'd138674130 :
   (i==6'd47) ? 30'd141688785 :
   (i==6'd48) ? 30'd144703440 :
   (i==6'd49) ? 30'd147718095 :
   (i==6'd50) ? 30'd150732750 :
   (i==6'd51) ? 30'd153747405 :
   (i==6'd52) ? 30'd156762060 :
   (i==6'd53) ? 30'd159776715 :
   (i==6'd54) ? 30'd162791370 :
   (i==6'd55) ? 30'd165806025 :
   (i==6'd56) ? 30'd168820680 :
   (i==6'd57) ? 30'd171835335 :
   (i==6'd58) ? 30'd174849990 :
   (i==6'd59) ? 30'd177864645 :
   (i==6'd60) ? 30'd180879300 :
   (i==6'd61) ? 30'd183893955 :
   (i==6'd62) ? 30'd186908610 :
   30'd189923265;

endmodule

module reduction_table_q1071513601(i, table_out);
input [5:0] i;
output [29:0] table_out;
assign table_out = 
   (i==6'd0) ? 30'd0 :
   (i==6'd1) ? 30'd2228223 :
   (i==6'd2) ? 30'd4456446 :
   (i==6'd3) ? 30'd6684669 :
   (i==6'd4) ? 30'd8912892 :
   (i==6'd5) ? 30'd11141115 :
   (i==6'd6) ? 30'd13369338 :
   (i==6'd7) ? 30'd15597561 :
   (i==6'd8) ? 30'd17825784 :
   (i==6'd9) ? 30'd20054007 :
   (i==6'd10) ? 30'd22282230 :
   (i==6'd11) ? 30'd24510453 :
   (i==6'd12) ? 30'd26738676 :
   (i==6'd13) ? 30'd28966899 :
   (i==6'd14) ? 30'd31195122 :
   (i==6'd15) ? 30'd33423345 :
   (i==6'd16) ? 30'd35651568 :
   (i==6'd17) ? 30'd37879791 :
   (i==6'd18) ? 30'd40108014 :
   (i==6'd19) ? 30'd42336237 :
   (i==6'd20) ? 30'd44564460 :
   (i==6'd21) ? 30'd46792683 :
   (i==6'd22) ? 30'd49020906 :
   (i==6'd23) ? 30'd51249129 :
   (i==6'd24) ? 30'd53477352 :
   (i==6'd25) ? 30'd55705575 :
   (i==6'd26) ? 30'd57933798 :
   (i==6'd27) ? 30'd60162021 :
   (i==6'd28) ? 30'd62390244 :
   (i==6'd29) ? 30'd64618467 :
   (i==6'd30) ? 30'd66846690 :
   (i==6'd31) ? 30'd69074913 :
   (i==6'd32) ? 30'd71303136 :
   (i==6'd33) ? 30'd73531359 :
   (i==6'd34) ? 30'd75759582 :
   (i==6'd35) ? 30'd77987805 :
   (i==6'd36) ? 30'd80216028 :
   (i==6'd37) ? 30'd82444251 :
   (i==6'd38) ? 30'd84672474 :
   (i==6'd39) ? 30'd86900697 :
   (i==6'd40) ? 30'd89128920 :
   (i==6'd41) ? 30'd91357143 :
   (i==6'd42) ? 30'd93585366 :
   (i==6'd43) ? 30'd95813589 :
   (i==6'd44) ? 30'd98041812 :
   (i==6'd45) ? 30'd100270035 :
   (i==6'd46) ? 30'd102498258 :
   (i==6'd47) ? 30'd104726481 :
   (i==6'd48) ? 30'd106954704 :
   (i==6'd49) ? 30'd109182927 :
   (i==6'd50) ? 30'd111411150 :
   (i==6'd51) ? 30'd113639373 :
   (i==6'd52) ? 30'd115867596 :
   (i==6'd53) ? 30'd118095819 :
   (i==6'd54) ? 30'd120324042 :
   (i==6'd55) ? 30'd122552265 :
   (i==6'd56) ? 30'd124780488 :
   (i==6'd57) ? 30'd127008711 :
   (i==6'd58) ? 30'd129236934 :
   (i==6'd59) ? 30'd131465157 :
   (i==6'd60) ? 30'd133693380 :
   (i==6'd61) ? 30'd135921603 :
   (i==6'd62) ? 30'd138149826 :
   30'd140378049;

endmodule

module reduction_table_q1072496641(i, table_out);
input [5:0] i;
output [29:0] table_out;
assign table_out = 
   (i==6'd0) ? 30'd0 :
   (i==6'd1) ? 30'd1245183 :
   (i==6'd2) ? 30'd2490366 :
   (i==6'd3) ? 30'd3735549 :
   (i==6'd4) ? 30'd4980732 :
   (i==6'd5) ? 30'd6225915 :
   (i==6'd6) ? 30'd7471098 :
   (i==6'd7) ? 30'd8716281 :
   (i==6'd8) ? 30'd9961464 :
   (i==6'd9) ? 30'd11206647 :
   (i==6'd10) ? 30'd12451830 :
   (i==6'd11) ? 30'd13697013 :
   (i==6'd12) ? 30'd14942196 :
   (i==6'd13) ? 30'd16187379 :
   (i==6'd14) ? 30'd17432562 :
   (i==6'd15) ? 30'd18677745 :
   (i==6'd16) ? 30'd19922928 :
   (i==6'd17) ? 30'd21168111 :
   (i==6'd18) ? 30'd22413294 :
   (i==6'd19) ? 30'd23658477 :
   (i==6'd20) ? 30'd24903660 :
   (i==6'd21) ? 30'd26148843 :
   (i==6'd22) ? 30'd27394026 :
   (i==6'd23) ? 30'd28639209 :
   (i==6'd24) ? 30'd29884392 :
   (i==6'd25) ? 30'd31129575 :
   (i==6'd26) ? 30'd32374758 :
   (i==6'd27) ? 30'd33619941 :
   (i==6'd28) ? 30'd34865124 :
   (i==6'd29) ? 30'd36110307 :
   (i==6'd30) ? 30'd37355490 :
   (i==6'd31) ? 30'd38600673 :
   (i==6'd32) ? 30'd39845856 :
   (i==6'd33) ? 30'd41091039 :
   (i==6'd34) ? 30'd42336222 :
   (i==6'd35) ? 30'd43581405 :
   (i==6'd36) ? 30'd44826588 :
   (i==6'd37) ? 30'd46071771 :
   (i==6'd38) ? 30'd47316954 :
   (i==6'd39) ? 30'd48562137 :
   (i==6'd40) ? 30'd49807320 :
   (i==6'd41) ? 30'd51052503 :
   (i==6'd42) ? 30'd52297686 :
   (i==6'd43) ? 30'd53542869 :
   (i==6'd44) ? 30'd54788052 :
   (i==6'd45) ? 30'd56033235 :
   (i==6'd46) ? 30'd57278418 :
   (i==6'd47) ? 30'd58523601 :
   (i==6'd48) ? 30'd59768784 :
   (i==6'd49) ? 30'd61013967 :
   (i==6'd50) ? 30'd62259150 :
   (i==6'd51) ? 30'd63504333 :
   (i==6'd52) ? 30'd64749516 :
   (i==6'd53) ? 30'd65994699 :
   (i==6'd54) ? 30'd67239882 :
   (i==6'd55) ? 30'd68485065 :
   (i==6'd56) ? 30'd69730248 :
   (i==6'd57) ? 30'd70975431 :
   (i==6'd58) ? 30'd72220614 :
   (i==6'd59) ? 30'd73465797 :
   (i==6'd60) ? 30'd74710980 :
   (i==6'd61) ? 30'd75956163 :
   (i==6'd62) ? 30'd77201346 :
   30'd78446529;

endmodule

module reduction_table_q1073479681(i, table_out);
input [5:0] i;
output [29:0] table_out;
assign table_out = 
   (i==6'd0) ? 30'd0 :
   (i==6'd1) ? 30'd262143 :
   (i==6'd2) ? 30'd524286 :
   (i==6'd3) ? 30'd786429 :
   (i==6'd4) ? 30'd1048572 :
   (i==6'd5) ? 30'd1310715 :
   (i==6'd6) ? 30'd1572858 :
   (i==6'd7) ? 30'd1835001 :
   (i==6'd8) ? 30'd2097144 :
   (i==6'd9) ? 30'd2359287 :
   (i==6'd10) ? 30'd2621430 :
   (i==6'd11) ? 30'd2883573 :
   (i==6'd12) ? 30'd3145716 :
   (i==6'd13) ? 30'd3407859 :
   (i==6'd14) ? 30'd3670002 :
   (i==6'd15) ? 30'd3932145 :
   (i==6'd16) ? 30'd4194288 :
   (i==6'd17) ? 30'd4456431 :
   (i==6'd18) ? 30'd4718574 :
   (i==6'd19) ? 30'd4980717 :
   (i==6'd20) ? 30'd5242860 :
   (i==6'd21) ? 30'd5505003 :
   (i==6'd22) ? 30'd5767146 :
   (i==6'd23) ? 30'd6029289 :
   (i==6'd24) ? 30'd6291432 :
   (i==6'd25) ? 30'd6553575 :
   (i==6'd26) ? 30'd6815718 :
   (i==6'd27) ? 30'd7077861 :
   (i==6'd28) ? 30'd7340004 :
   (i==6'd29) ? 30'd7602147 :
   (i==6'd30) ? 30'd7864290 :
   (i==6'd31) ? 30'd8126433 :
   (i==6'd32) ? 30'd8388576 :
   (i==6'd33) ? 30'd8650719 :
   (i==6'd34) ? 30'd8912862 :
   (i==6'd35) ? 30'd9175005 :
   (i==6'd36) ? 30'd9437148 :
   (i==6'd37) ? 30'd9699291 :
   (i==6'd38) ? 30'd9961434 :
   (i==6'd39) ? 30'd10223577 :
   (i==6'd40) ? 30'd10485720 :
   (i==6'd41) ? 30'd10747863 :
   (i==6'd42) ? 30'd11010006 :
   (i==6'd43) ? 30'd11272149 :
   (i==6'd44) ? 30'd11534292 :
   (i==6'd45) ? 30'd11796435 :
   (i==6'd46) ? 30'd12058578 :
   (i==6'd47) ? 30'd12320721 :
   (i==6'd48) ? 30'd12582864 :
   (i==6'd49) ? 30'd12845007 :
   (i==6'd50) ? 30'd13107150 :
   (i==6'd51) ? 30'd13369293 :
   (i==6'd52) ? 30'd13631436 :
   (i==6'd53) ? 30'd13893579 :
   (i==6'd54) ? 30'd14155722 :
   (i==6'd55) ? 30'd14417865 :
   (i==6'd56) ? 30'd14680008 :
   (i==6'd57) ? 30'd14942151 :
   (i==6'd58) ? 30'd15204294 :
   (i==6'd59) ? 30'd15466437 :
   (i==6'd60) ? 30'd15728580 :
   (i==6'd61) ? 30'd15990723 :
   (i==6'd62) ? 30'd16252866 :
   30'd16515009;

endmodule

module reduction_table_q1068433409(i, table_out);
input [5:0] i;
output [29:0] table_out;
assign table_out = 
   (i==6'd0) ? 30'd0 :
   (i==6'd1) ? 30'd5308415 :
   (i==6'd2) ? 30'd10616830 :
   (i==6'd3) ? 30'd15925245 :
   (i==6'd4) ? 30'd21233660 :
   (i==6'd5) ? 30'd26542075 :
   (i==6'd6) ? 30'd31850490 :
   (i==6'd7) ? 30'd37158905 :
   (i==6'd8) ? 30'd42467320 :
   (i==6'd9) ? 30'd47775735 :
   (i==6'd10) ? 30'd53084150 :
   (i==6'd11) ? 30'd58392565 :
   (i==6'd12) ? 30'd63700980 :
   (i==6'd13) ? 30'd69009395 :
   (i==6'd14) ? 30'd74317810 :
   (i==6'd15) ? 30'd79626225 :
   (i==6'd16) ? 30'd84934640 :
   (i==6'd17) ? 30'd90243055 :
   (i==6'd18) ? 30'd95551470 :
   (i==6'd19) ? 30'd100859885 :
   (i==6'd20) ? 30'd106168300 :
   (i==6'd21) ? 30'd111476715 :
   (i==6'd22) ? 30'd116785130 :
   (i==6'd23) ? 30'd122093545 :
   (i==6'd24) ? 30'd127401960 :
   (i==6'd25) ? 30'd132710375 :
   (i==6'd26) ? 30'd138018790 :
   (i==6'd27) ? 30'd143327205 :
   (i==6'd28) ? 30'd148635620 :
   (i==6'd29) ? 30'd153944035 :
   (i==6'd30) ? 30'd159252450 :
   (i==6'd31) ? 30'd164560865 :
   (i==6'd32) ? 30'd169869280 :
   (i==6'd33) ? 30'd175177695 :
   (i==6'd34) ? 30'd180486110 :
   (i==6'd35) ? 30'd185794525 :
   (i==6'd36) ? 30'd191102940 :
   (i==6'd37) ? 30'd196411355 :
   (i==6'd38) ? 30'd201719770 :
   (i==6'd39) ? 30'd207028185 :
   (i==6'd40) ? 30'd212336600 :
   (i==6'd41) ? 30'd217645015 :
   (i==6'd42) ? 30'd222953430 :
   (i==6'd43) ? 30'd228261845 :
   (i==6'd44) ? 30'd233570260 :
   (i==6'd45) ? 30'd238878675 :
   (i==6'd46) ? 30'd244187090 :
   (i==6'd47) ? 30'd249495505 :
   (i==6'd48) ? 30'd254803920 :
   (i==6'd49) ? 30'd260112335 :
   (i==6'd50) ? 30'd265420750 :
   (i==6'd51) ? 30'd270729165 :
   (i==6'd52) ? 30'd276037580 :
   (i==6'd53) ? 30'd281345995 :
   (i==6'd54) ? 30'd286654410 :
   (i==6'd55) ? 30'd291962825 :
   (i==6'd56) ? 30'd297271240 :
   (i==6'd57) ? 30'd302579655 :
   (i==6'd58) ? 30'd307888070 :
   (i==6'd59) ? 30'd313196485 :
   (i==6'd60) ? 30'd318504900 :
   (i==6'd61) ? 30'd323813315 :
   (i==6'd62) ? 30'd329121730 :
   30'd334430145;

endmodule

module reduction_table_q1068236801(i, table_out);
input [5:0] i;
output [29:0] table_out;
assign table_out = 
   (i==6'd0) ? 30'd0 :
   (i==6'd1) ? 30'd5505023 :
   (i==6'd2) ? 30'd11010046 :
   (i==6'd3) ? 30'd16515069 :
   (i==6'd4) ? 30'd22020092 :
   (i==6'd5) ? 30'd27525115 :
   (i==6'd6) ? 30'd33030138 :
   (i==6'd7) ? 30'd38535161 :
   (i==6'd8) ? 30'd44040184 :
   (i==6'd9) ? 30'd49545207 :
   (i==6'd10) ? 30'd55050230 :
   (i==6'd11) ? 30'd60555253 :
   (i==6'd12) ? 30'd66060276 :
   (i==6'd13) ? 30'd71565299 :
   (i==6'd14) ? 30'd77070322 :
   (i==6'd15) ? 30'd82575345 :
   (i==6'd16) ? 30'd88080368 :
   (i==6'd17) ? 30'd93585391 :
   (i==6'd18) ? 30'd99090414 :
   (i==6'd19) ? 30'd104595437 :
   (i==6'd20) ? 30'd110100460 :
   (i==6'd21) ? 30'd115605483 :
   (i==6'd22) ? 30'd121110506 :
   (i==6'd23) ? 30'd126615529 :
   (i==6'd24) ? 30'd132120552 :
   (i==6'd25) ? 30'd137625575 :
   (i==6'd26) ? 30'd143130598 :
   (i==6'd27) ? 30'd148635621 :
   (i==6'd28) ? 30'd154140644 :
   (i==6'd29) ? 30'd159645667 :
   (i==6'd30) ? 30'd165150690 :
   (i==6'd31) ? 30'd170655713 :
   (i==6'd32) ? 30'd176160736 :
   (i==6'd33) ? 30'd181665759 :
   (i==6'd34) ? 30'd187170782 :
   (i==6'd35) ? 30'd192675805 :
   (i==6'd36) ? 30'd198180828 :
   (i==6'd37) ? 30'd203685851 :
   (i==6'd38) ? 30'd209190874 :
   (i==6'd39) ? 30'd214695897 :
   (i==6'd40) ? 30'd220200920 :
   (i==6'd41) ? 30'd225705943 :
   (i==6'd42) ? 30'd231210966 :
   (i==6'd43) ? 30'd236715989 :
   (i==6'd44) ? 30'd242221012 :
   (i==6'd45) ? 30'd247726035 :
   (i==6'd46) ? 30'd253231058 :
   (i==6'd47) ? 30'd258736081 :
   (i==6'd48) ? 30'd264241104 :
   (i==6'd49) ? 30'd269746127 :
   (i==6'd50) ? 30'd275251150 :
   (i==6'd51) ? 30'd280756173 :
   (i==6'd52) ? 30'd286261196 :
   (i==6'd53) ? 30'd291766219 :
   (i==6'd54) ? 30'd297271242 :
   (i==6'd55) ? 30'd302776265 :
   (i==6'd56) ? 30'd308281288 :
   (i==6'd57) ? 30'd313786311 :
   (i==6'd58) ? 30'd319291334 :
   (i==6'd59) ? 30'd324796357 :
   (i==6'd60) ? 30'd330301380 :
   (i==6'd61) ? 30'd335806403 :
   (i==6'd62) ? 30'd341311426 :
   30'd346816449;

endmodule

module reduction_table_q1065811969(i, table_out);
input [5:0] i;
output [29:0] table_out;
assign table_out = 
   (i==6'd0) ? 30'd0 :
   (i==6'd1) ? 30'd7929855 :
   (i==6'd2) ? 30'd15859710 :
   (i==6'd3) ? 30'd23789565 :
   (i==6'd4) ? 30'd31719420 :
   (i==6'd5) ? 30'd39649275 :
   (i==6'd6) ? 30'd47579130 :
   (i==6'd7) ? 30'd55508985 :
   (i==6'd8) ? 30'd63438840 :
   (i==6'd9) ? 30'd71368695 :
   (i==6'd10) ? 30'd79298550 :
   (i==6'd11) ? 30'd87228405 :
   (i==6'd12) ? 30'd95158260 :
   (i==6'd13) ? 30'd103088115 :
   (i==6'd14) ? 30'd111017970 :
   (i==6'd15) ? 30'd118947825 :
   (i==6'd16) ? 30'd126877680 :
   (i==6'd17) ? 30'd134807535 :
   (i==6'd18) ? 30'd142737390 :
   (i==6'd19) ? 30'd150667245 :
   (i==6'd20) ? 30'd158597100 :
   (i==6'd21) ? 30'd166526955 :
   (i==6'd22) ? 30'd174456810 :
   (i==6'd23) ? 30'd182386665 :
   (i==6'd24) ? 30'd190316520 :
   (i==6'd25) ? 30'd198246375 :
   (i==6'd26) ? 30'd206176230 :
   (i==6'd27) ? 30'd214106085 :
   (i==6'd28) ? 30'd222035940 :
   (i==6'd29) ? 30'd229965795 :
   (i==6'd30) ? 30'd237895650 :
   (i==6'd31) ? 30'd245825505 :
   (i==6'd32) ? 30'd253755360 :
   (i==6'd33) ? 30'd261685215 :
   (i==6'd34) ? 30'd269615070 :
   (i==6'd35) ? 30'd277544925 :
   (i==6'd36) ? 30'd285474780 :
   (i==6'd37) ? 30'd293404635 :
   (i==6'd38) ? 30'd301334490 :
   (i==6'd39) ? 30'd309264345 :
   (i==6'd40) ? 30'd317194200 :
   (i==6'd41) ? 30'd325124055 :
   (i==6'd42) ? 30'd333053910 :
   (i==6'd43) ? 30'd340983765 :
   (i==6'd44) ? 30'd348913620 :
   (i==6'd45) ? 30'd356843475 :
   (i==6'd46) ? 30'd364773330 :
   (i==6'd47) ? 30'd372703185 :
   (i==6'd48) ? 30'd380633040 :
   (i==6'd49) ? 30'd388562895 :
   (i==6'd50) ? 30'd396492750 :
   (i==6'd51) ? 30'd404422605 :
   (i==6'd52) ? 30'd412352460 :
   (i==6'd53) ? 30'd420282315 :
   (i==6'd54) ? 30'd428212170 :
   (i==6'd55) ? 30'd436142025 :
   (i==6'd56) ? 30'd444071880 :
   (i==6'd57) ? 30'd452001735 :
   (i==6'd58) ? 30'd459931590 :
   (i==6'd59) ? 30'd467861445 :
   (i==6'd60) ? 30'd475791300 :
   (i==6'd61) ? 30'd483721155 :
   (i==6'd62) ? 30'd491651010 :
   30'd499580865;

endmodule

module reduction_table_q1065484289(i, table_out);
input [5:0] i;
output [29:0] table_out;
assign table_out = 
   (i==6'd0) ? 30'd0 :
   (i==6'd1) ? 30'd8257535 :
   (i==6'd2) ? 30'd16515070 :
   (i==6'd3) ? 30'd24772605 :
   (i==6'd4) ? 30'd33030140 :
   (i==6'd5) ? 30'd41287675 :
   (i==6'd6) ? 30'd49545210 :
   (i==6'd7) ? 30'd57802745 :
   (i==6'd8) ? 30'd66060280 :
   (i==6'd9) ? 30'd74317815 :
   (i==6'd10) ? 30'd82575350 :
   (i==6'd11) ? 30'd90832885 :
   (i==6'd12) ? 30'd99090420 :
   (i==6'd13) ? 30'd107347955 :
   (i==6'd14) ? 30'd115605490 :
   (i==6'd15) ? 30'd123863025 :
   (i==6'd16) ? 30'd132120560 :
   (i==6'd17) ? 30'd140378095 :
   (i==6'd18) ? 30'd148635630 :
   (i==6'd19) ? 30'd156893165 :
   (i==6'd20) ? 30'd165150700 :
   (i==6'd21) ? 30'd173408235 :
   (i==6'd22) ? 30'd181665770 :
   (i==6'd23) ? 30'd189923305 :
   (i==6'd24) ? 30'd198180840 :
   (i==6'd25) ? 30'd206438375 :
   (i==6'd26) ? 30'd214695910 :
   (i==6'd27) ? 30'd222953445 :
   (i==6'd28) ? 30'd231210980 :
   (i==6'd29) ? 30'd239468515 :
   (i==6'd30) ? 30'd247726050 :
   (i==6'd31) ? 30'd255983585 :
   (i==6'd32) ? 30'd264241120 :
   (i==6'd33) ? 30'd272498655 :
   (i==6'd34) ? 30'd280756190 :
   (i==6'd35) ? 30'd289013725 :
   (i==6'd36) ? 30'd297271260 :
   (i==6'd37) ? 30'd305528795 :
   (i==6'd38) ? 30'd313786330 :
   (i==6'd39) ? 30'd322043865 :
   (i==6'd40) ? 30'd330301400 :
   (i==6'd41) ? 30'd338558935 :
   (i==6'd42) ? 30'd346816470 :
   (i==6'd43) ? 30'd355074005 :
   (i==6'd44) ? 30'd363331540 :
   (i==6'd45) ? 30'd371589075 :
   (i==6'd46) ? 30'd379846610 :
   (i==6'd47) ? 30'd388104145 :
   (i==6'd48) ? 30'd396361680 :
   (i==6'd49) ? 30'd404619215 :
   (i==6'd50) ? 30'd412876750 :
   (i==6'd51) ? 30'd421134285 :
   (i==6'd52) ? 30'd429391820 :
   (i==6'd53) ? 30'd437649355 :
   (i==6'd54) ? 30'd445906890 :
   (i==6'd55) ? 30'd454164425 :
   (i==6'd56) ? 30'd462421960 :
   (i==6'd57) ? 30'd470679495 :
   (i==6'd58) ? 30'd478937030 :
   (i==6'd59) ? 30'd487194565 :
   (i==6'd60) ? 30'd495452100 :
   (i==6'd61) ? 30'd503709635 :
   (i==6'd62) ? 30'd511967170 :
   30'd520224705;

endmodule

module reduction_table_q1064697857(i, table_out);
input [5:0] i;
output [29:0] table_out;
assign table_out = 
   (i==6'd0) ? 30'd0 :
   (i==6'd1) ? 30'd9043967 :
   (i==6'd2) ? 30'd18087934 :
   (i==6'd3) ? 30'd27131901 :
   (i==6'd4) ? 30'd36175868 :
   (i==6'd5) ? 30'd45219835 :
   (i==6'd6) ? 30'd54263802 :
   (i==6'd7) ? 30'd63307769 :
   (i==6'd8) ? 30'd72351736 :
   (i==6'd9) ? 30'd81395703 :
   (i==6'd10) ? 30'd90439670 :
   (i==6'd11) ? 30'd99483637 :
   (i==6'd12) ? 30'd108527604 :
   (i==6'd13) ? 30'd117571571 :
   (i==6'd14) ? 30'd126615538 :
   (i==6'd15) ? 30'd135659505 :
   (i==6'd16) ? 30'd144703472 :
   (i==6'd17) ? 30'd153747439 :
   (i==6'd18) ? 30'd162791406 :
   (i==6'd19) ? 30'd171835373 :
   (i==6'd20) ? 30'd180879340 :
   (i==6'd21) ? 30'd189923307 :
   (i==6'd22) ? 30'd198967274 :
   (i==6'd23) ? 30'd208011241 :
   (i==6'd24) ? 30'd217055208 :
   (i==6'd25) ? 30'd226099175 :
   (i==6'd26) ? 30'd235143142 :
   (i==6'd27) ? 30'd244187109 :
   (i==6'd28) ? 30'd253231076 :
   (i==6'd29) ? 30'd262275043 :
   (i==6'd30) ? 30'd271319010 :
   (i==6'd31) ? 30'd280362977 :
   (i==6'd32) ? 30'd289406944 :
   (i==6'd33) ? 30'd298450911 :
   (i==6'd34) ? 30'd307494878 :
   (i==6'd35) ? 30'd316538845 :
   (i==6'd36) ? 30'd325582812 :
   (i==6'd37) ? 30'd334626779 :
   (i==6'd38) ? 30'd343670746 :
   (i==6'd39) ? 30'd352714713 :
   (i==6'd40) ? 30'd361758680 :
   (i==6'd41) ? 30'd370802647 :
   (i==6'd42) ? 30'd379846614 :
   (i==6'd43) ? 30'd388890581 :
   (i==6'd44) ? 30'd397934548 :
   (i==6'd45) ? 30'd406978515 :
   (i==6'd46) ? 30'd416022482 :
   (i==6'd47) ? 30'd425066449 :
   (i==6'd48) ? 30'd434110416 :
   (i==6'd49) ? 30'd443154383 :
   (i==6'd50) ? 30'd452198350 :
   (i==6'd51) ? 30'd461242317 :
   (i==6'd52) ? 30'd470286284 :
   (i==6'd53) ? 30'd479330251 :
   (i==6'd54) ? 30'd488374218 :
   (i==6'd55) ? 30'd497418185 :
   (i==6'd56) ? 30'd506462152 :
   (i==6'd57) ? 30'd515506119 :
   (i==6'd58) ? 30'd524550086 :
   (i==6'd59) ? 30'd533594053 :
   (i==6'd60) ? 30'd542638020 :
   (i==6'd61) ? 30'd551681987 :
   (i==6'd62) ? 30'd560725954 :
   30'd569769921;

endmodule

module reduction_table_q1063452673(i, table_out);
input [5:0] i;
output [29:0] table_out;
assign table_out = 
   (i==6'd0) ? 30'd0 :
   (i==6'd1) ? 30'd10289151 :
   (i==6'd2) ? 30'd20578302 :
   (i==6'd3) ? 30'd30867453 :
   (i==6'd4) ? 30'd41156604 :
   (i==6'd5) ? 30'd51445755 :
   (i==6'd6) ? 30'd61734906 :
   (i==6'd7) ? 30'd72024057 :
   (i==6'd8) ? 30'd82313208 :
   (i==6'd9) ? 30'd92602359 :
   (i==6'd10) ? 30'd102891510 :
   (i==6'd11) ? 30'd113180661 :
   (i==6'd12) ? 30'd123469812 :
   (i==6'd13) ? 30'd133758963 :
   (i==6'd14) ? 30'd144048114 :
   (i==6'd15) ? 30'd154337265 :
   (i==6'd16) ? 30'd164626416 :
   (i==6'd17) ? 30'd174915567 :
   (i==6'd18) ? 30'd185204718 :
   (i==6'd19) ? 30'd195493869 :
   (i==6'd20) ? 30'd205783020 :
   (i==6'd21) ? 30'd216072171 :
   (i==6'd22) ? 30'd226361322 :
   (i==6'd23) ? 30'd236650473 :
   (i==6'd24) ? 30'd246939624 :
   (i==6'd25) ? 30'd257228775 :
   (i==6'd26) ? 30'd267517926 :
   (i==6'd27) ? 30'd277807077 :
   (i==6'd28) ? 30'd288096228 :
   (i==6'd29) ? 30'd298385379 :
   (i==6'd30) ? 30'd308674530 :
   (i==6'd31) ? 30'd318963681 :
   (i==6'd32) ? 30'd329252832 :
   (i==6'd33) ? 30'd339541983 :
   (i==6'd34) ? 30'd349831134 :
   (i==6'd35) ? 30'd360120285 :
   (i==6'd36) ? 30'd370409436 :
   (i==6'd37) ? 30'd380698587 :
   (i==6'd38) ? 30'd390987738 :
   (i==6'd39) ? 30'd401276889 :
   (i==6'd40) ? 30'd411566040 :
   (i==6'd41) ? 30'd421855191 :
   (i==6'd42) ? 30'd432144342 :
   (i==6'd43) ? 30'd442433493 :
   (i==6'd44) ? 30'd452722644 :
   (i==6'd45) ? 30'd463011795 :
   (i==6'd46) ? 30'd473300946 :
   (i==6'd47) ? 30'd483590097 :
   (i==6'd48) ? 30'd493879248 :
   (i==6'd49) ? 30'd504168399 :
   (i==6'd50) ? 30'd514457550 :
   (i==6'd51) ? 30'd524746701 :
   (i==6'd52) ? 30'd535035852 :
   (i==6'd53) ? 30'd545325003 :
   (i==6'd54) ? 30'd555614154 :
   (i==6'd55) ? 30'd565903305 :
   (i==6'd56) ? 30'd576192456 :
   (i==6'd57) ? 30'd586481607 :
   (i==6'd58) ? 30'd596770758 :
   (i==6'd59) ? 30'd607059909 :
   (i==6'd60) ? 30'd617349060 :
   (i==6'd61) ? 30'd627638211 :
   (i==6'd62) ? 30'd637927362 :
   30'd648216513;

endmodule


module reduction_table_q1063321601(i, table_out);
input [5:0] i;
output [29:0] table_out;
assign table_out = 
   (i==6'd0) ? 30'd0 :
   (i==6'd1) ? 30'd10420223 :
   (i==6'd2) ? 30'd20840446 :
   (i==6'd3) ? 30'd31260669 :
   (i==6'd4) ? 30'd41680892 :
   (i==6'd5) ? 30'd52101115 :
   (i==6'd6) ? 30'd62521338 :
   (i==6'd7) ? 30'd72941561 :
   (i==6'd8) ? 30'd83361784 :
   (i==6'd9) ? 30'd93782007 :
   (i==6'd10) ? 30'd104202230 :
   (i==6'd11) ? 30'd114622453 :
   (i==6'd12) ? 30'd125042676 :
   (i==6'd13) ? 30'd135462899 :
   (i==6'd14) ? 30'd145883122 :
   (i==6'd15) ? 30'd156303345 :
   (i==6'd16) ? 30'd166723568 :
   (i==6'd17) ? 30'd177143791 :
   (i==6'd18) ? 30'd187564014 :
   (i==6'd19) ? 30'd197984237 :
   (i==6'd20) ? 30'd208404460 :
   (i==6'd21) ? 30'd218824683 :
   (i==6'd22) ? 30'd229244906 :
   (i==6'd23) ? 30'd239665129 :
   (i==6'd24) ? 30'd250085352 :
   (i==6'd25) ? 30'd260505575 :
   (i==6'd26) ? 30'd270925798 :
   (i==6'd27) ? 30'd281346021 :
   (i==6'd28) ? 30'd291766244 :
   (i==6'd29) ? 30'd302186467 :
   (i==6'd30) ? 30'd312606690 :
   (i==6'd31) ? 30'd323026913 :
   (i==6'd32) ? 30'd333447136 :
   (i==6'd33) ? 30'd343867359 :
   (i==6'd34) ? 30'd354287582 :
   (i==6'd35) ? 30'd364707805 :
   (i==6'd36) ? 30'd375128028 :
   (i==6'd37) ? 30'd385548251 :
   (i==6'd38) ? 30'd395968474 :
   (i==6'd39) ? 30'd406388697 :
   (i==6'd40) ? 30'd416808920 :
   (i==6'd41) ? 30'd427229143 :
   (i==6'd42) ? 30'd437649366 :
   (i==6'd43) ? 30'd448069589 :
   (i==6'd44) ? 30'd458489812 :
   (i==6'd45) ? 30'd468910035 :
   (i==6'd46) ? 30'd479330258 :
   (i==6'd47) ? 30'd489750481 :
   (i==6'd48) ? 30'd500170704 :
   (i==6'd49) ? 30'd510590927 :
   (i==6'd50) ? 30'd521011150 :
   (i==6'd51) ? 30'd531431373 :
   (i==6'd52) ? 30'd541851596 :
   (i==6'd53) ? 30'd552271819 :
   (i==6'd54) ? 30'd562692042 :
   (i==6'd55) ? 30'd573112265 :
   (i==6'd56) ? 30'd583532488 :
   (i==6'd57) ? 30'd593952711 :
   (i==6'd58) ? 30'd604372934 :
   (i==6'd59) ? 30'd614793157 :
   (i==6'd60) ? 30'd625213380 :
   (i==6'd61) ? 30'd635633603 :
   (i==6'd62) ? 30'd646053826 :
   30'd656474049;

endmodule

